`timescale 1ns / 1ps
// Calculations are performed using fixed-point representation,
// with 2 integer bits and WIDTH-2 fractional bits,
// formatted as xx.xxxxxx
module psi #(
    parameter WIDTH = 8  // Bit Width should be between 5 and 8
) (
    input  wire [WIDTH-1:0] psi_in,
    output reg  [WIDTH-1:0] psi_out
);

  always @(psi_in) begin
    case (WIDTH)
      5: begin
        case (psi_in)
          5'b00000: psi_out <= 5'b11111;
          5'b00001: psi_out <= 5'b10110;
          5'b00010: psi_out <= 5'b10001;
          5'b00011: psi_out <= 5'b01101;
          5'b00100: psi_out <= 5'b01011;
          5'b00101: psi_out <= 5'b01010;
          5'b00110: psi_out <= 5'b01000;
          5'b00111: psi_out <= 5'b00111;
          5'b01000: psi_out <= 5'b00110;
          5'b01001: psi_out <= 5'b00101;
          5'b01010: psi_out <= 5'b00101;
          5'b01011: psi_out <= 5'b00100;
          5'b01100: psi_out <= 5'b00100;
          5'b01101: psi_out <= 5'b00011;
          5'b01110: psi_out <= 5'b00011;
          5'b01111: psi_out <= 5'b00010;
          5'b10000: psi_out <= 5'b00010;
          5'b10001: psi_out <= 5'b00010;
          5'b10010: psi_out <= 5'b00010;
          5'b10011: psi_out <= 5'b00001;
          5'b10100: psi_out <= 5'b00001;
          5'b10101: psi_out <= 5'b00001;
          5'b10110: psi_out <= 5'b00001;
          5'b10111: psi_out <= 5'b00001;
          5'b11000: psi_out <= 5'b00001;
          5'b11001: psi_out <= 5'b00001;
          5'b11010: psi_out <= 5'b00001;
          5'b11011: psi_out <= 5'b00001;
          5'b11100: psi_out <= 5'b00000;
          5'b11101: psi_out <= 5'b00000;
          5'b11110: psi_out <= 5'b00000;
          5'b11111: psi_out <= 5'b00000;
          // default:  psi_out <= 5'b00000;
        endcase
      end
      6: begin
        case (psi_in)
          6'b000000: psi_out <= 6'b111111;
          6'b000001: psi_out <= 6'b110111;
          6'b000010: psi_out <= 6'b101100;
          6'b000011: psi_out <= 6'b100110;
          6'b000100: psi_out <= 6'b100001;
          6'b000101: psi_out <= 6'b011110;
          6'b000110: psi_out <= 6'b011011;
          6'b000111: psi_out <= 6'b011001;
          6'b001000: psi_out <= 6'b010111;
          6'b001001: psi_out <= 6'b010101;
          6'b001010: psi_out <= 6'b010011;
          6'b001011: psi_out <= 6'b010010;
          6'b001100: psi_out <= 6'b010000;
          6'b001101: psi_out <= 6'b001111;
          6'b001110: psi_out <= 6'b001110;
          6'b001111: psi_out <= 6'b001101;
          6'b010000: psi_out <= 6'b001100;
          6'b010001: psi_out <= 6'b001100;
          6'b010010: psi_out <= 6'b001011;
          6'b010011: psi_out <= 6'b001010;
          6'b010100: psi_out <= 6'b001001;
          6'b010101: psi_out <= 6'b001001;
          6'b010110: psi_out <= 6'b001000;
          6'b010111: psi_out <= 6'b001000;
          6'b011000: psi_out <= 6'b000111;
          6'b011001: psi_out <= 6'b000111;
          6'b011010: psi_out <= 6'b000110;
          6'b011011: psi_out <= 6'b000110;
          6'b011100: psi_out <= 6'b000110;
          6'b011101: psi_out <= 6'b000101;
          6'b011110: psi_out <= 6'b000101;
          6'b011111: psi_out <= 6'b000101;
          6'b100000: psi_out <= 6'b000100;
          6'b100001: psi_out <= 6'b000100;
          6'b100010: psi_out <= 6'b000100;
          6'b100011: psi_out <= 6'b000100;
          6'b100100: psi_out <= 6'b000011;
          6'b100101: psi_out <= 6'b000011;
          6'b100110: psi_out <= 6'b000011;
          6'b100111: psi_out <= 6'b000011;
          6'b101000: psi_out <= 6'b000011;
          6'b101001: psi_out <= 6'b000010;
          6'b101010: psi_out <= 6'b000010;
          6'b101011: psi_out <= 6'b000010;
          6'b101100: psi_out <= 6'b000010;
          6'b101101: psi_out <= 6'b000010;
          6'b101110: psi_out <= 6'b000010;
          6'b101111: psi_out <= 6'b000010;
          6'b110000: psi_out <= 6'b000010;
          6'b110001: psi_out <= 6'b000001;
          6'b110010: psi_out <= 6'b000001;
          6'b110011: psi_out <= 6'b000001;
          6'b110100: psi_out <= 6'b000001;
          6'b110101: psi_out <= 6'b000001;
          6'b110110: psi_out <= 6'b000001;
          6'b110111: psi_out <= 6'b000001;
          6'b111000: psi_out <= 6'b000001;
          6'b111001: psi_out <= 6'b000001;
          6'b111010: psi_out <= 6'b000001;
          6'b111011: psi_out <= 6'b000001;
          6'b111100: psi_out <= 6'b000001;
          6'b111101: psi_out <= 6'b000001;
          6'b111110: psi_out <= 6'b000001;
          6'b111111: psi_out <= 6'b000000;
          // default:   psi_out <= 6'b000000;
        endcase
      end
      // 7: begin
      //   case (psi_in)
      //     7'b0000000: psi_out <= 7'b1111111;
      //     7'b0000001: psi_out <= 7'b1111111;
      //     7'b0000010: psi_out <= 7'b1101111;
      //     7'b0000011: psi_out <= 7'b1100010;
      //     7'b0000100: psi_out <= 7'b1011001;
      //     7'b0000101: psi_out <= 7'b1010010;
      //     7'b0000110: psi_out <= 7'b1001100;
      //     7'b0000111: psi_out <= 7'b1000111;
      //     7'b0001000: psi_out <= 7'b1000011;
      //     7'b0001001: psi_out <= 7'b0111111;
      //     7'b0001010: psi_out <= 7'b0111100;
      //     7'b0001011: psi_out <= 7'b0111001;
      //     7'b0001100: psi_out <= 7'b0110110;
      //     7'b0001101: psi_out <= 7'b0110011;
      //     7'b0001110: psi_out <= 7'b0110001;
      //     7'b0001111: psi_out <= 7'b0101111;
      //     7'b0010000: psi_out <= 7'b0101101;
      //     7'b0010001: psi_out <= 7'b0101011;
      //     7'b0010010: psi_out <= 7'b0101001;
      //     7'b0010011: psi_out <= 7'b0101000;
      //     7'b0010100: psi_out <= 7'b0100110;
      //     7'b0010101: psi_out <= 7'b0100101;
      //     7'b0010110: psi_out <= 7'b0100011;
      //     7'b0010111: psi_out <= 7'b0100010;
      //     7'b0011000: psi_out <= 7'b0100001;
      //     7'b0011001: psi_out <= 7'b0100000;
      //     7'b0011010: psi_out <= 7'b0011111;
      //     7'b0011011: psi_out <= 7'b0011101;
      //     7'b0011100: psi_out <= 7'b0011100;
      //     7'b0011101: psi_out <= 7'b0011011;
      //     7'b0011110: psi_out <= 7'b0011010;
      //     7'b0011111: psi_out <= 7'b0011010;
      //     7'b0100000: psi_out <= 7'b0011001;
      //     7'b0100001: psi_out <= 7'b0011000;
      //     7'b0100010: psi_out <= 7'b0010111;
      //     7'b0100011: psi_out <= 7'b0010110;
      //     7'b0100100: psi_out <= 7'b0010110;
      //     7'b0100101: psi_out <= 7'b0010101;
      //     7'b0100110: psi_out <= 7'b0010100;
      //     7'b0100111: psi_out <= 7'b0010100;
      //     7'b0101000: psi_out <= 7'b0010011;
      //     7'b0101001: psi_out <= 7'b0010010;
      //     7'b0101010: psi_out <= 7'b0010010;
      //     7'b0101011: psi_out <= 7'b0010001;
      //     7'b0101100: psi_out <= 7'b0010001;
      //     7'b0101101: psi_out <= 7'b0010000;
      //     7'b0101110: psi_out <= 7'b0001111;
      //     7'b0101111: psi_out <= 7'b0001111;
      //     7'b0110000: psi_out <= 7'b0001111;
      //     7'b0110001: psi_out <= 7'b0001110;
      //     7'b0110010: psi_out <= 7'b0001110;
      //     7'b0110011: psi_out <= 7'b0001101;
      //     7'b0110100: psi_out <= 7'b0001101;
      //     7'b0110101: psi_out <= 7'b0001100;
      //     7'b0110110: psi_out <= 7'b0001100;
      //     7'b0110111: psi_out <= 7'b0001100;
      //     7'b0111000: psi_out <= 7'b0001011;
      //     7'b0111001: psi_out <= 7'b0001011;
      //     7'b0111010: psi_out <= 7'b0001011;
      //     7'b0111011: psi_out <= 7'b0001010;
      //     7'b0111100: psi_out <= 7'b0001010;
      //     7'b0111101: psi_out <= 7'b0001010;
      //     7'b0111110: psi_out <= 7'b0001001;
      //     7'b0111111: psi_out <= 7'b0001001;
      //     7'b1000000: psi_out <= 7'b0001001;
      //     7'b1000001: psi_out <= 7'b0001000;
      //     7'b1000010: psi_out <= 7'b0001000;
      //     7'b1000011: psi_out <= 7'b0001000;
      //     7'b1000100: psi_out <= 7'b0001000;
      //     7'b1000101: psi_out <= 7'b0000111;
      //     7'b1000110: psi_out <= 7'b0000111;
      //     7'b1000111: psi_out <= 7'b0000111;
      //     7'b1001000: psi_out <= 7'b0000111;
      //     7'b1001001: psi_out <= 7'b0000111;
      //     7'b1001010: psi_out <= 7'b0000110;
      //     7'b1001011: psi_out <= 7'b0000110;
      //     7'b1001100: psi_out <= 7'b0000110;
      //     7'b1001101: psi_out <= 7'b0000110;
      //     7'b1001110: psi_out <= 7'b0000110;
      //     7'b1001111: psi_out <= 7'b0000101;
      //     7'b1010000: psi_out <= 7'b0000101;
      //     7'b1010001: psi_out <= 7'b0000101;
      //     7'b1010010: psi_out <= 7'b0000101;
      //     7'b1010011: psi_out <= 7'b0000101;
      //     7'b1010100: psi_out <= 7'b0000101;
      //     7'b1010101: psi_out <= 7'b0000101;
      //     7'b1010110: psi_out <= 7'b0000100;
      //     7'b1010111: psi_out <= 7'b0000100;
      //     7'b1011000: psi_out <= 7'b0000100;
      //     7'b1011001: psi_out <= 7'b0000100;
      //     7'b1011010: psi_out <= 7'b0000100;
      //     7'b1011011: psi_out <= 7'b0000100;
      //     7'b1011100: psi_out <= 7'b0000100;
      //     7'b1011101: psi_out <= 7'b0000100;
      //     7'b1011110: psi_out <= 7'b0000011;
      //     7'b1011111: psi_out <= 7'b0000011;
      //     7'b1100000: psi_out <= 7'b0000011;
      //     7'b1100001: psi_out <= 7'b0000011;
      //     7'b1100010: psi_out <= 7'b0000011;
      //     7'b1100011: psi_out <= 7'b0000011;
      //     7'b1100100: psi_out <= 7'b0000011;
      //     7'b1100101: psi_out <= 7'b0000011;
      //     7'b1100110: psi_out <= 7'b0000011;
      //     7'b1100111: psi_out <= 7'b0000011;
      //     7'b1101000: psi_out <= 7'b0000010;
      //     7'b1101001: psi_out <= 7'b0000010;
      //     7'b1101010: psi_out <= 7'b0000010;
      //     7'b1101011: psi_out <= 7'b0000010;
      //     7'b1101100: psi_out <= 7'b0000010;
      //     7'b1101101: psi_out <= 7'b0000010;
      //     7'b1101110: psi_out <= 7'b0000010;
      //     7'b1101111: psi_out <= 7'b0000010;
      //     7'b1110000: psi_out <= 7'b0000010;
      //     7'b1110001: psi_out <= 7'b0000010;
      //     7'b1110010: psi_out <= 7'b0000010;
      //     7'b1110011: psi_out <= 7'b0000010;
      //     7'b1110100: psi_out <= 7'b0000010;
      //     7'b1110101: psi_out <= 7'b0000010;
      //     7'b1110110: psi_out <= 7'b0000010;
      //     7'b1110111: psi_out <= 7'b0000010;
      //     7'b1111000: psi_out <= 7'b0000010;
      //     7'b1111001: psi_out <= 7'b0000001;
      //     7'b1111010: psi_out <= 7'b0000001;
      //     7'b1111011: psi_out <= 7'b0000001;
      //     7'b1111100: psi_out <= 7'b0000001;
      //     7'b1111101: psi_out <= 7'b0000001;
      //     7'b1111110: psi_out <= 7'b0000001;
      //     7'b1111111: psi_out <= 7'b0000000;
      //     default: psi_out <= 7'b0000000;
      //   endcase
      // end
      // 8: begin
      //   case (psi_in)
      //     8'b00000000: psi_out <= 8'b11111111;
      //     8'b00000001: psi_out <= 8'b11111111;
      //     8'b00000010: psi_out <= 8'b11111111;
      //     8'b00000011: psi_out <= 8'b11110000;
      //     8'b00000100: psi_out <= 8'b11011110;
      //     8'b00000101: psi_out <= 8'b11010000;
      //     8'b00000110: psi_out <= 8'b11000100;
      //     8'b00000111: psi_out <= 8'b10111010;
      //     8'b00001000: psi_out <= 8'b10110010;
      //     8'b00001001: psi_out <= 8'b10101010;
      //     8'b00001010: psi_out <= 8'b10100011;
      //     8'b00001011: psi_out <= 8'b10011101;
      //     8'b00001100: psi_out <= 8'b10011000;
      //     8'b00001101: psi_out <= 8'b10010011;
      //     8'b00001110: psi_out <= 8'b10001110;
      //     8'b00001111: psi_out <= 8'b10001010;
      //     8'b00010000: psi_out <= 8'b10000101;
      //     8'b00010001: psi_out <= 8'b10000010;
      //     8'b00010010: psi_out <= 8'b01111110;
      //     8'b00010011: psi_out <= 8'b01111011;
      //     8'b00010100: psi_out <= 8'b01110111;
      //     8'b00010101: psi_out <= 8'b01110100;
      //     8'b00010110: psi_out <= 8'b01110001;
      //     8'b00010111: psi_out <= 8'b01101111;
      //     8'b00011000: psi_out <= 8'b01101100;
      //     8'b00011001: psi_out <= 8'b01101001;
      //     8'b00011010: psi_out <= 8'b01100111;
      //     8'b00011011: psi_out <= 8'b01100101;
      //     8'b00011100: psi_out <= 8'b01100010;
      //     8'b00011101: psi_out <= 8'b01100000;
      //     8'b00011110: psi_out <= 8'b01011110;
      //     8'b00011111: psi_out <= 8'b01011100;
      //     8'b00100000: psi_out <= 8'b01011010;
      //     8'b00100001: psi_out <= 8'b01011000;
      //     8'b00100010: psi_out <= 8'b01010110;
      //     8'b00100011: psi_out <= 8'b01010101;
      //     8'b00100100: psi_out <= 8'b01010011;
      //     8'b00100101: psi_out <= 8'b01010001;
      //     8'b00100110: psi_out <= 8'b01010000;
      //     8'b00100111: psi_out <= 8'b01001110;
      //     8'b00101000: psi_out <= 8'b01001100;
      //     8'b00101001: psi_out <= 8'b01001011;
      //     8'b00101010: psi_out <= 8'b01001010;
      //     8'b00101011: psi_out <= 8'b01001000;
      //     8'b00101100: psi_out <= 8'b01000111;
      //     8'b00101101: psi_out <= 8'b01000101;
      //     8'b00101110: psi_out <= 8'b01000100;
      //     8'b00101111: psi_out <= 8'b01000011;
      //     8'b00110000: psi_out <= 8'b01000010;
      //     8'b00110001: psi_out <= 8'b01000000;
      //     8'b00110010: psi_out <= 8'b00111111;
      //     8'b00110011: psi_out <= 8'b00111110;
      //     8'b00110100: psi_out <= 8'b00111101;
      //     8'b00110101: psi_out <= 8'b00111100;
      //     8'b00110110: psi_out <= 8'b00111011;
      //     8'b00110111: psi_out <= 8'b00111010;
      //     8'b00111000: psi_out <= 8'b00111001;
      //     8'b00111001: psi_out <= 8'b00111000;
      //     8'b00111010: psi_out <= 8'b00110111;
      //     8'b00111011: psi_out <= 8'b00110110;
      //     8'b00111100: psi_out <= 8'b00110101;
      //     8'b00111101: psi_out <= 8'b00110100;
      //     8'b00111110: psi_out <= 8'b00110011;
      //     8'b00111111: psi_out <= 8'b00110010;
      //     8'b01000000: psi_out <= 8'b00110001;
      //     8'b01000001: psi_out <= 8'b00110001;
      //     8'b01000010: psi_out <= 8'b00110000;
      //     8'b01000011: psi_out <= 8'b00101111;
      //     8'b01000100: psi_out <= 8'b00101110;
      //     8'b01000101: psi_out <= 8'b00101101;
      //     8'b01000110: psi_out <= 8'b00101101;
      //     8'b01000111: psi_out <= 8'b00101100;
      //     8'b01001000: psi_out <= 8'b00101011;
      //     8'b01001001: psi_out <= 8'b00101010;
      //     8'b01001010: psi_out <= 8'b00101010;
      //     8'b01001011: psi_out <= 8'b00101001;
      //     8'b01001100: psi_out <= 8'b00101000;
      //     8'b01001101: psi_out <= 8'b00101000;
      //     8'b01001110: psi_out <= 8'b00100111;
      //     8'b01001111: psi_out <= 8'b00100110;
      //     8'b01010000: psi_out <= 8'b00100110;
      //     8'b01010001: psi_out <= 8'b00100101;
      //     8'b01010010: psi_out <= 8'b00100101;
      //     8'b01010011: psi_out <= 8'b00100100;
      //     8'b01010100: psi_out <= 8'b00100011;
      //     8'b01010101: psi_out <= 8'b00100011;
      //     8'b01010110: psi_out <= 8'b00100010;
      //     8'b01010111: psi_out <= 8'b00100010;
      //     8'b01011000: psi_out <= 8'b00100001;
      //     8'b01011001: psi_out <= 8'b00100001;
      //     8'b01011010: psi_out <= 8'b00100000;
      //     8'b01011011: psi_out <= 8'b00100000;
      //     8'b01011100: psi_out <= 8'b00011111;
      //     8'b01011101: psi_out <= 8'b00011110;
      //     8'b01011110: psi_out <= 8'b00011110;
      //     8'b01011111: psi_out <= 8'b00011110;
      //     8'b01100000: psi_out <= 8'b00011101;
      //     8'b01100001: psi_out <= 8'b00011101;
      //     8'b01100010: psi_out <= 8'b00011100;
      //     8'b01100011: psi_out <= 8'b00011100;
      //     8'b01100100: psi_out <= 8'b00011011;
      //     8'b01100101: psi_out <= 8'b00011011;
      //     8'b01100110: psi_out <= 8'b00011010;
      //     8'b01100111: psi_out <= 8'b00011010;
      //     8'b01101000: psi_out <= 8'b00011010;
      //     8'b01101001: psi_out <= 8'b00011001;
      //     8'b01101010: psi_out <= 8'b00011001;
      //     8'b01101011: psi_out <= 8'b00011000;
      //     8'b01101100: psi_out <= 8'b00011000;
      //     8'b01101101: psi_out <= 8'b00011000;
      //     8'b01101110: psi_out <= 8'b00010111;
      //     8'b01101111: psi_out <= 8'b00010111;
      //     8'b01110000: psi_out <= 8'b00010110;
      //     8'b01110001: psi_out <= 8'b00010110;
      //     8'b01110010: psi_out <= 8'b00010110;
      //     8'b01110011: psi_out <= 8'b00010101;
      //     8'b01110100: psi_out <= 8'b00010101;
      //     8'b01110101: psi_out <= 8'b00010101;
      //     8'b01110110: psi_out <= 8'b00010100;
      //     8'b01110111: psi_out <= 8'b00010100;
      //     8'b01111000: psi_out <= 8'b00010100;
      //     8'b01111001: psi_out <= 8'b00010011;
      //     8'b01111010: psi_out <= 8'b00010011;
      //     8'b01111011: psi_out <= 8'b00010011;
      //     8'b01111100: psi_out <= 8'b00010011;
      //     8'b01111101: psi_out <= 8'b00010010;
      //     8'b01111110: psi_out <= 8'b00010010;
      //     8'b01111111: psi_out <= 8'b00010010;
      //     8'b10000000: psi_out <= 8'b00010001;
      //     8'b10000001: psi_out <= 8'b00010001;
      //     8'b10000010: psi_out <= 8'b00010001;
      //     8'b10000011: psi_out <= 8'b00010001;
      //     8'b10000100: psi_out <= 8'b00010000;
      //     8'b10000101: psi_out <= 8'b00010000;
      //     8'b10000110: psi_out <= 8'b00010000;
      //     8'b10000111: psi_out <= 8'b00010000;
      //     8'b10001000: psi_out <= 8'b00001111;
      //     8'b10001001: psi_out <= 8'b00001111;
      //     8'b10001010: psi_out <= 8'b00001111;
      //     8'b10001011: psi_out <= 8'b00001111;
      //     8'b10001100: psi_out <= 8'b00001110;
      //     8'b10001101: psi_out <= 8'b00001110;
      //     8'b10001110: psi_out <= 8'b00001110;
      //     8'b10001111: psi_out <= 8'b00001110;
      //     8'b10010000: psi_out <= 8'b00001110;
      //     8'b10010001: psi_out <= 8'b00001101;
      //     8'b10010010: psi_out <= 8'b00001101;
      //     8'b10010011: psi_out <= 8'b00001101;
      //     8'b10010100: psi_out <= 8'b00001101;
      //     8'b10010101: psi_out <= 8'b00001101;
      //     8'b10010110: psi_out <= 8'b00001100;
      //     8'b10010111: psi_out <= 8'b00001100;
      //     8'b10011000: psi_out <= 8'b00001100;
      //     8'b10011001: psi_out <= 8'b00001100;
      //     8'b10011010: psi_out <= 8'b00001100;
      //     8'b10011011: psi_out <= 8'b00001011;
      //     8'b10011100: psi_out <= 8'b00001011;
      //     8'b10011101: psi_out <= 8'b00001011;
      //     8'b10011110: psi_out <= 8'b00001011;
      //     8'b10011111: psi_out <= 8'b00001011;
      //     8'b10100000: psi_out <= 8'b00001011;
      //     8'b10100001: psi_out <= 8'b00001010;
      //     8'b10100010: psi_out <= 8'b00001010;
      //     8'b10100011: psi_out <= 8'b00001010;
      //     8'b10100100: psi_out <= 8'b00001010;
      //     8'b10100101: psi_out <= 8'b00001010;
      //     8'b10100110: psi_out <= 8'b00001010;
      //     8'b10100111: psi_out <= 8'b00001001;
      //     8'b10101000: psi_out <= 8'b00001001;
      //     8'b10101001: psi_out <= 8'b00001001;
      //     8'b10101010: psi_out <= 8'b00001001;
      //     8'b10101011: psi_out <= 8'b00001001;
      //     8'b10101100: psi_out <= 8'b00001001;
      //     8'b10101101: psi_out <= 8'b00001001;
      //     8'b10101110: psi_out <= 8'b00001000;
      //     8'b10101111: psi_out <= 8'b00001000;
      //     8'b10110000: psi_out <= 8'b00001000;
      //     8'b10110001: psi_out <= 8'b00001000;
      //     8'b10110010: psi_out <= 8'b00001000;
      //     8'b10110011: psi_out <= 8'b00001000;
      //     8'b10110100: psi_out <= 8'b00001000;
      //     8'b10110101: psi_out <= 8'b00001000;
      //     8'b10110110: psi_out <= 8'b00000111;
      //     8'b10110111: psi_out <= 8'b00000111;
      //     8'b10111000: psi_out <= 8'b00000111;
      //     8'b10111001: psi_out <= 8'b00000111;
      //     8'b10111010: psi_out <= 8'b00000111;
      //     8'b10111011: psi_out <= 8'b00000111;
      //     8'b10111100: psi_out <= 8'b00000111;
      //     8'b10111101: psi_out <= 8'b00000111;
      //     8'b10111110: psi_out <= 8'b00000111;
      //     8'b10111111: psi_out <= 8'b00000110;
      //     8'b11000000: psi_out <= 8'b00000110;
      //     8'b11000001: psi_out <= 8'b00000110;
      //     8'b11000010: psi_out <= 8'b00000110;
      //     8'b11000011: psi_out <= 8'b00000110;
      //     8'b11000100: psi_out <= 8'b00000110;
      //     8'b11000101: psi_out <= 8'b00000110;
      //     8'b11000110: psi_out <= 8'b00000110;
      //     8'b11000111: psi_out <= 8'b00000110;
      //     8'b11001000: psi_out <= 8'b00000110;
      //     8'b11001001: psi_out <= 8'b00000110;
      //     8'b11001010: psi_out <= 8'b00000101;
      //     8'b11001011: psi_out <= 8'b00000101;
      //     8'b11001100: psi_out <= 8'b00000101;
      //     8'b11001101: psi_out <= 8'b00000101;
      //     8'b11001110: psi_out <= 8'b00000101;
      //     8'b11001111: psi_out <= 8'b00000101;
      //     8'b11010000: psi_out <= 8'b00000101;
      //     8'b11010001: psi_out <= 8'b00000101;
      //     8'b11010010: psi_out <= 8'b00000101;
      //     8'b11010011: psi_out <= 8'b00000101;
      //     8'b11010100: psi_out <= 8'b00000101;
      //     8'b11010101: psi_out <= 8'b00000101;
      //     8'b11010110: psi_out <= 8'b00000101;
      //     8'b11010111: psi_out <= 8'b00000100;
      //     8'b11011000: psi_out <= 8'b00000100;
      //     8'b11011001: psi_out <= 8'b00000100;
      //     8'b11011010: psi_out <= 8'b00000100;
      //     8'b11011011: psi_out <= 8'b00000100;
      //     8'b11011100: psi_out <= 8'b00000100;
      //     8'b11011101: psi_out <= 8'b00000100;
      //     8'b11011110: psi_out <= 8'b00000100;
      //     8'b11011111: psi_out <= 8'b00000100;
      //     8'b11100000: psi_out <= 8'b00000100;
      //     8'b11100001: psi_out <= 8'b00000100;
      //     8'b11100010: psi_out <= 8'b00000100;
      //     8'b11100011: psi_out <= 8'b00000100;
      //     8'b11100100: psi_out <= 8'b00000100;
      //     8'b11100101: psi_out <= 8'b00000100;
      //     8'b11100110: psi_out <= 8'b00000100;
      //     8'b11100111: psi_out <= 8'b00000011;
      //     8'b11101000: psi_out <= 8'b00000011;
      //     8'b11101001: psi_out <= 8'b00000011;
      //     8'b11101010: psi_out <= 8'b00000011;
      //     8'b11101011: psi_out <= 8'b00000011;
      //     8'b11101100: psi_out <= 8'b00000011;
      //     8'b11101101: psi_out <= 8'b00000011;
      //     8'b11101110: psi_out <= 8'b00000011;
      //     8'b11101111: psi_out <= 8'b00000011;
      //     8'b11110000: psi_out <= 8'b00000011;
      //     8'b11110001: psi_out <= 8'b00000011;
      //     8'b11110010: psi_out <= 8'b00000011;
      //     8'b11110011: psi_out <= 8'b00000011;
      //     8'b11110100: psi_out <= 8'b00000011;
      //     8'b11110101: psi_out <= 8'b00000011;
      //     8'b11110110: psi_out <= 8'b00000011;
      //     8'b11110111: psi_out <= 8'b00000011;
      //     8'b11111000: psi_out <= 8'b00000011;
      //     8'b11111001: psi_out <= 8'b00000011;
      //     8'b11111010: psi_out <= 8'b00000011;
      //     8'b11111011: psi_out <= 8'b00000011;
      //     8'b11111100: psi_out <= 8'b00000010;
      //     8'b11111101: psi_out <= 8'b00000010;
      //     8'b11111110: psi_out <= 8'b00000010;
      //     8'b11111111: psi_out <= 8'b00000000;
      //     default: psi_out <= 8'b00000000;
      //   endcase
      // end
    endcase
  end
endmodule
