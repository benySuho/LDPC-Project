`timescale 1ns / 1ps
`define INPUT_FILE "../input/matrix.txt"

module ldpc_decoder_tb;

  // Parameters
  parameter MAX_BLOCK_SIZE = 64;
  parameter MAX_ROWS = 12;
  parameter MAX_COLS = 24;
  parameter MAX_ITERATIONS = 50;
  parameter WIDTH_LLR = 6;
  parameter INITIAL_LLR = 5'b10110;
  localparam MAX_CODE_LEN = MAX_COLS * MAX_BLOCK_SIZE;
  localparam MAX_MSG_LEN = MAX_ROWS * MAX_BLOCK_SIZE;
  localparam WIDTH_CODE_LEN = $clog2(MAX_CODE_LEN + 1);
  localparam WIDTH_BLOCK = $clog2(MAX_BLOCK_SIZE);
  localparam WIDTH_ROWS = $clog2(MAX_ROWS + 1);
  localparam WIDTH_COLS = $clog2(MAX_COLS + 1);
  localparam WIDTH_ITERATION = $clog2(MAX_ITERATIONS + 1);

  // Inputs
  reg clk;
  reg rst_n;
  reg start_conf_input;
  reg start_input;
  // reg [WIDTH_CODE_LEN-1:0] codeword_len_in;
  reg [MAX_CODE_LEN-1:0] codeword_in;
  reg [MAX_CODE_LEN-1:0] original;
  reg [MAX_CODE_LEN-1:0] codeword_out;
  reg [MAX_CODE_LEN-1:0] codeword_inital;
  reg [MAX_ROWS*MAX_COLS*WIDTH_BLOCK-1:0] h_matrix_in;
  reg [WIDTH_BLOCK-1:0] block_size_in;
  reg [WIDTH_ROWS-1:0] rows_in;
  reg [WIDTH_COLS-1:0] cols_in;
  reg [WIDTH_ITERATION-1:0] iterations_in;
  reg [MAX_BLOCK_SIZE-1:0] data_in, data_out;
  reg [MAX_BLOCK_SIZE-1:0] temp_num;

  // Outputs
  wire [MAX_CODE_LEN-1:0] estimate;
  wire valid;
  wire done;

  integer i, j, i_max;
  integer data_file;
  integer scan_file;
  integer num;

  // Instantiate the DUT (Device Under Test)
  ldpc_decoder #(
      .MAX_BLOCK_SIZE(MAX_BLOCK_SIZE),
      .MAX_ROWS(MAX_ROWS),
      .MAX_COLS(MAX_COLS),
      .MAX_ITERATIONS(MAX_ITERATIONS),
      .WIDTH_LLR(WIDTH_LLR),
      .INITIAL_LLR(INITIAL_LLR)
  ) decoder (
      .clk(clk),
      .rst_n(rst_n),
      .start_input(start_input),
      .start_conf_input(start_conf_input),
      .data_in(data_in),
      .data_out(data_out),
      .valid(valid),
      .done(done)
  );

  // Clock generation
  initial begin
    clk = 1;
    forever #5 clk = ~clk;  // 10 ns clock period
  end

  // Test stimulus
  initial begin
    // Initialize inputs
    rst_n = 0;
    // codeword_len_in = 0;
    codeword_in = 0;
    original = 0;
    codeword_inital = 0;
    h_matrix_in = 0;
    block_size_in = 0;
    rows_in = 0;
    cols_in = 0;
    iterations_in = 0;
    start_conf_input = 0;
    start_input = 0;

    // Apply reset
    #10 rst_n = 1;


    data_file = $fopen(`INPUT_FILE, "r");
    if (data_file == 0) begin
      $display("Error: Could not open file.");
      $finish;
    end


    scan_file = $fscanf(data_file, "%d\n", num);
    rows_in = num;
    scan_file = $fscanf(data_file, "%d\n", num);
    cols_in = num;
    scan_file = $fscanf(data_file, "%d\n", num);
    block_size_in = num;

    // input matrix
    h_matrix_in = {(MAX_COLS * MAX_COLS * WIDTH_BLOCK) {1'b1}};

    for (i = 0; i < rows_in; i++) begin
      for (j = 0; j < cols_in; j++) begin
        scan_file = $fscanf(data_file, "%d\n", num);
        if (num == -1) begin
          h_matrix_in[(i*MAX_COLS+j)*WIDTH_BLOCK+:WIDTH_BLOCK] = {(WIDTH_BLOCK) {1'b1}};
        end else begin
          h_matrix_in[(i*MAX_COLS+j)*WIDTH_BLOCK+:WIDTH_BLOCK] = num % MAX_BLOCK_SIZE;
        end
      end
    end

    $display("Rows: %d, Columns: %d, Block Size: %d", rows_in, cols_in, block_size_in);

    $fclose(data_file);

    iterations_in = 50;  // Maximum iterations (50)

    data_in = 0;
    data_in[7:0] = {(8) {1'b0}} | rows_in;
    data_in[15:8] = {(8) {1'b0}} | cols_in;
    data_in[23:16] = {(8) {1'b0}} | iterations_in;
    data_in[31:24] = {(8) {1'b0}} | block_size_in;
    start_conf_input = 1;
    #10 start_conf_input = 0;
    #20;
    i_max = ((MAX_COLS * MAX_ROWS * WIDTH_BLOCK + MAX_BLOCK_SIZE - 1) / MAX_BLOCK_SIZE);
    for (i = 0; i < i_max; i = i + 1) begin
      if (i == i_max - 1) begin
        start_conf_input = 1;
        data_in = h_matrix_in[MAX_COLS*MAX_ROWS*WIDTH_BLOCK-1:MAX_COLS*MAX_ROWS*WIDTH_BLOCK-1-MAX_BLOCK_SIZE];
      end else begin
        data_in = {(MAX_BLOCK_SIZE) {1'b0}} | h_matrix_in[i*MAX_BLOCK_SIZE+:MAX_BLOCK_SIZE];
      end
      #10;
    end

    start_conf_input = 0;

    $display("1: Expected Success");
    // input codeword
    original = 1368'b101111100010000001111011011111110001111110001000111110101110011101111010100010100111001110001110111100101100100000110001101001000010111001010111110100101110100010000110001110011001111101000000111000111100000011001010001011101101000111100001011000111010111101111100000111010101101101010011110110100000000101111011111100100111011011000110001001101111010000010000100001011000010010010101001101110101001110101111111111101001101100011011100001111011100111000101010000111001000100111100001100110000110000111110100010001111000010000011001100001110001100000101110110001111100000101111101100001100100101100011011110100101011101110000010101100101100101111011100001011000111101111100000000000001110000010011011100010110010010010011111000111011010111111010010100001110001010111010100100111001100100000010011101101011100010001010010100101110010000111111001110010001000110110100101101001101111110110111000000100001011110100010100111101110001111010010000001000100000111110110010001001111000111101111000100100111101111001011000010011110100111101110011100111011110110101111001110110011100010101000000100101101011011010101110011001110001001010010110110011101101100101101101110000101010010010011111110010111101101101000000101100101110101000110010110000110111110101100011011101111110010001101010001111100000101000110100110101111010011110100101110001000011010101100011000111010110100101011;
    codeword_in = 1368'b101011100010000001111011111111110001111110001000111110101110011101101010100010100111001110001110110100111100100000110001101001000010101001010111110100101110100010000110101110011001111101000000111000111100000011001010001011101101000101100001011000111010111101111100001111010101101101010011110111100000000101111011111100100111011011100110001001101111010000010000110001011000010010010101001101110101001110101111111111101001101100011011110001111011100111000101010000111001000100111100001100110000110000111110100010001111000010000011001100001110001100000101110110001111100000101111101100001100100101100011011110100101011101110000010101000101101101111011100001011000111101111100000000000001110000010011011100010110010010010011111000111011010111111010010100001110101110111010100100111001100100000010011100101011100010000010010100101110010000111111001110010001000110110100001101001101110110110111000000000001011110100010100111101110001111010010000001000100000111110110010011001111000111101111000100100111101111001011000011011110100111101110011100111011110110101111001110110001100010101000000110101101011011010101110011001110001001010010110110011001101100101101100110000101010010010001111110011111101101101000000101100101110101000110010110000110111110101100011011101111110010001101010001111100000101000110100010101111010011110100101110001000011010101100011000111010110100001011;
    // $display("5: Expected Fail");
    // // input codeword
    // original = 1368'b101000111011100010111111000010010011011100100001110010000001111001001110101011110100111111010011001111010100000101111110110011000010101010001010100011010110011011011101110110000011100101010001110110010000100110010110101001110111101101100001011111000001001101110000110011110011000011111101001000001100000101111110101111010011110000100111011000111001011100001111011100100111100010000001000101101011000111010001100011101011100011100100111011101001001010010111000000101100011111101000111100011010110100111101110111001111001001111011101011101101111000010011110100001001111110010110111111011111011101010001111011011000100011100000011010111010011111011000000001010111111100000101001100100000111100001011011011001010100111011010111110010010111001000101101101001000011010111000010111101001100001101100001010100001101000001010110010011110001110000001000101111010101001010010110010101011100111001101111010001100101101001110111100101100010010011001010000111010110010010101100111101110110101110000111001010010001101011100010110011011111000000001010011000100000110100111101100000110101011100010110101100100111110101110111010010100010001101010010111111010010110011000010100011100110010100100010010011010110111110010101011111011011100111001010100010000100101001001000110110101010111000011010011101010000001110001111011111100010000111101111011100000101011110010011101011110111000001001;
    // codeword_in = 1368'b101001111011100010111111000010010011011100100001110010000001111001001110101011110100111111010011001110010100000101111110110011000010101010001010100011010110111011011101110110000011100101010001110110010000100110010110101101110111101101100001011111000001001101110000110011110011000011111101001001001100000101101110101111010011110000100110011000111001011100001111011100100111100010000001000101101011000111010001100011101011100011100100011011101001001010010111000000101000011111101000111100011010110100111101110111001111001001111011101011101001111000010111110100001001100110010110111111001111011101010001111011011000100011110000011010111010011111011000000001010111111101000101001000100000011000001011111011001010100111011010111110010110111001000101101001001000011010111000010111101001100001101100001010100001101000001010110010011110001110000000000101111010101000010010110010101011100111001101111010001100101101001100111100101100010010011001010000111010110010010001100111101110110101110000111001010011001101011100010110011011111000001001010011000100000110100111101100100110101011100010110101100100111110101111111010010100010001101010010111110010000110011000010100011000110010100100010010011010110111110010100011111011011100111001110101010000100101001001000110110101010111000011010011101000000000110000111011111100010000111101111011100000111011110010011101011110111000001001;

    // Process decode
    send_codeword(codeword_in);
    wait (done);
    receive_codeword();
    print_result();


    // Stop simulation
    #100 $finish;
  end

  task automatic send_codeword;
    input [MAX_COLS*MAX_BLOCK_SIZE-1:0] codeword;  // Input codeword

    integer i;  // Loop variable
    reg [MAX_BLOCK_SIZE-1:0] temp_num;

    begin
      #10 start_input = 1;
      #10 start_input = 0;
      #10;
      for (i = 0; i < MAX_COLS; i = i + 1) begin
        if (i < cols_in) begin
          temp_num = codeword[MAX_BLOCK_SIZE-1:0];
          temp_num = temp_num << (MAX_BLOCK_SIZE - block_size_in);
          codeword = codeword >> block_size_in;
          data_in  = temp_num;
        end else begin
          data_in = 0;
        end
        #10;  // Simulation delay
      end
    end
  endtask

  task automatic receive_codeword;
    codeword_out = 0;
    for (i = 0; i < MAX_COLS; i = i + 1) begin
      #10;
      codeword_out[i*block_size_in+:MAX_BLOCK_SIZE] = (data_out >> (MAX_BLOCK_SIZE-block_size_in));
    end
  endtask

  task automatic print_result;
    // Print vectors
    $display("%h", original);
    $display("%h", codeword_out);

    if (valid) begin
      $display("\tDecoded output is valid");
      if (codeword_out == original) begin
        $display("\tCodeword restored");
      end else begin
        $display("\tCodeword not restored");
      end
    end else begin
      $display("\tDecoding failed");
    end
  endtask

endmodule
