`timescale 1ns / 1ps
`define INPUT_FILE "../input/matrix.txt"

module ldpc_tb;

  // Parameters
  parameter MAX_BLOCK_SIZE = 64;
  parameter MAX_ROWS = 12;
  parameter MAX_COLS = 24;
  parameter MAX_ITERATIONS = 50;
  parameter WIDTH_LLR = 6;
  parameter INITIAL_LLR = 5'b10110;
  localparam MAX_CODE_LEN = MAX_COLS * MAX_BLOCK_SIZE;
  localparam MAX_MSG_LEN = MAX_ROWS * MAX_BLOCK_SIZE;
  localparam WIDTH_CODE_LEN = $clog2(MAX_CODE_LEN + 1);
  localparam WIDTH_BLOCK = $clog2(MAX_BLOCK_SIZE);
  localparam WIDTH_ROWS = $clog2(MAX_ROWS + 1);
  localparam WIDTH_COLS = $clog2(MAX_COLS + 1);
  localparam WIDTH_ITERATION = $clog2(MAX_ITERATIONS + 1);


  // Inputs
  reg clk;
  reg rst_n;
  reg start_conf_input_enc, start_conf_input_dec;
  reg start_input_enc, start_input_dec;
  reg [MAX_CODE_LEN-1:0] msg;
  reg [MAX_ROWS*MAX_COLS*WIDTH_BLOCK-1:0] matrix_in;
  reg [WIDTH_ROWS-1:0] rows_in;
  reg [WIDTH_COLS-1:0] cols_in;
  reg [WIDTH_BLOCK-1:0] block_size;
  reg [MAX_BLOCK_SIZE-1:0] data_in_enc, data_out_enc;
  reg [MAX_BLOCK_SIZE-1:0] data_in_dec, data_out_dec;
  reg [WIDTH_ITERATION-1:0] iterations_in;

  // Outputs
  reg [MAX_CODE_LEN-1:0] codeword, err_codeword;
  reg [MAX_CODE_LEN-1:0] rec_msg;
  reg [MAX_CODE_LEN-1:0] original;

  wire done_enc, done_dec;

  integer i, j, i_max;
  integer scan_file, data_file;
  integer num;


  // Instantiate the Encoder
  ldpc_encoder #(
      .MAX_BLOCK_SIZE(MAX_BLOCK_SIZE),
      .MAX_ROWS(MAX_ROWS),
      .MAX_COLS(MAX_COLS)
  ) encoder (
      .clk(clk),
      .rst_n(rst_n),
      .start_input(start_input_enc),
      .start_conf_input(start_conf_input_enc),
      .data_in(data_in_enc),
      .data_out(data_out_enc),
      .done(done_enc)
  );

  // Instantiate the Decoder
  ldpc_decoder #(
      .MAX_BLOCK_SIZE(MAX_BLOCK_SIZE),
      .MAX_ROWS(MAX_ROWS),
      .MAX_COLS(MAX_COLS),
      .MAX_ITERATIONS(MAX_ITERATIONS),
      .WIDTH_LLR(WIDTH_LLR),
      .INITIAL_LLR(INITIAL_LLR)
  ) decoder (
      .clk(clk),
      .rst_n(rst_n),
      .start_input(start_input_dec),
      .start_conf_input(start_conf_input_dec),
      .data_in(data_in_dec),
      .data_out(data_out_dec),
      .valid(valid),
      .done(done_dec)
  );

  // Clock generation
  initial begin
    clk = 1;
    forever #5 clk = ~clk;  // Toggle clock every 5 time units
  end

  // Testbench process
  initial begin
    // Initialize inputs
    rst_n = 0;
    msg = 0;
    matrix_in = 0;
    block_size = 0;
    rows_in = 0;
    cols_in = 0;
    start_conf_input_enc = 0;
    start_conf_input_dec = 0;
    start_input_enc = 0;
    start_input_dec = 0;

    // Apply reset
    #10 rst_n = 1;


    data_file = $fopen(`INPUT_FILE, "r");
    if (data_file == 0) begin
      $display("Error: Could not open file.");
      $finish;
    end


    scan_file = $fscanf(data_file, "%d\n", num);
    rows_in = num;
    scan_file = $fscanf(data_file, "%d\n", num);
    cols_in = num;
    scan_file = $fscanf(data_file, "%d\n", num);
    block_size = num;

    // input matrix
    matrix_in = {(MAX_COLS * MAX_COLS * WIDTH_BLOCK) {1'b1}};

    for (i = 0; i < rows_in; i++) begin
      for (j = 0; j < cols_in; j++) begin
        scan_file = $fscanf(data_file, "%d\n", num);
        if (num == -1) begin
          matrix_in[(i*MAX_COLS+j)*WIDTH_BLOCK+:WIDTH_BLOCK] = {(WIDTH_BLOCK) {1'b1}};
        end else begin
          matrix_in[(i*MAX_COLS+j)*WIDTH_BLOCK+:WIDTH_BLOCK] = num % block_size;
        end
      end
    end

    $fclose(data_file);

    // Send matrix to encoder
    data_in_enc = 0;
    data_in_enc[7:0] = {(8) {1'b0}} | rows_in;
    data_in_enc[15:8] = {(8) {1'b0}} | cols_in;
    data_in_enc[23:16] = {(8) {1'b0}} | block_size;
    start_conf_input_enc = 1;
    #10 start_conf_input_enc = 0;
    #20;
    i_max = ((MAX_COLS * MAX_ROWS * WIDTH_BLOCK + MAX_BLOCK_SIZE - 1) / MAX_BLOCK_SIZE);
    for (i = 0; i < i_max; i = i + 1) begin
      if (i == i_max - 1) begin
        start_conf_input_enc = 1;
        data_in_enc = matrix_in[MAX_COLS*MAX_ROWS*WIDTH_BLOCK-1:MAX_COLS*MAX_ROWS*WIDTH_BLOCK-1-MAX_BLOCK_SIZE];
      end else begin
        data_in_enc = {(MAX_BLOCK_SIZE) {1'b0}} | matrix_in[i*MAX_BLOCK_SIZE+:MAX_BLOCK_SIZE];
      end
      #10;
    end
    start_conf_input_enc = 0;

    // Send matrix to Decoder
    iterations_in = 50;  // Maximum iterations (50)
    data_in_dec = 0;
    data_in_dec[7:0] = {(8) {1'b0}} | rows_in;
    data_in_dec[15:8] = {(8) {1'b0}} | cols_in;
    data_in_dec[23:16] = {(8) {1'b0}} | iterations_in;
    data_in_dec[31:24] = {(8) {1'b0}} | block_size;
    start_conf_input_dec = 1;
    #10 start_conf_input_dec = 0;
    #20;
    i_max = ((MAX_COLS * MAX_ROWS * WIDTH_BLOCK + MAX_BLOCK_SIZE - 1) / MAX_BLOCK_SIZE);
    for (i = 0; i < i_max; i = i + 1) begin
      if (i == i_max - 1) begin
        start_conf_input_dec = 1;
        data_in_dec = matrix_in[MAX_COLS*MAX_ROWS*WIDTH_BLOCK-1:MAX_COLS*MAX_ROWS*WIDTH_BLOCK-1-MAX_BLOCK_SIZE];
      end else begin
        data_in_dec = {(MAX_BLOCK_SIZE) {1'b0}} | matrix_in[i*MAX_BLOCK_SIZE+:MAX_BLOCK_SIZE];
      end
      #10;
    end
    start_conf_input_dec = 0;

    // Input the message to be encoded, and encoded message for comparison
    // $display("1: Expected Fail");
    // // input codeword
    // msg = 1368'b101110110110100000011110100111010110110011001100000010111101100101110100011110111000101110010101111111100001100011000001011101100101110000011101010011110111110010111110110110100100010010011001000001101000010101010110001111001011101111100110011111110010110001011110101111011000010000011001011100111111000011101101000011001101011001110000101111110111110100100100111000110001000000111100001011100010110011010110101011100110100111110001011010100001110110011100110111001101110100100111010101011001000000100101101000001100010000001000010010000110101001111011111101011111110010011001010011000000110110101011011110110111011111111001111001101100101010010011101000010101010011000000011000011000100000101101111100100110011010001111101010001101101010110001010011110101111001100100010101000100111001000011101011111111011100001000110000111010100111101001111000111010010110000111000100111011000100010000010110110111011000111001111000101111011010011100010010111010110100110110110111110110100001110110011001001010010100100011010100111000100111;
    // original = 1368'b101110110110100000011110100111010110110011001100000010111101100101110100011110111000101110010101111111100001100011000001011101100101110000011101010011110111110010111110110110100100010010011001000001101000010101010110001111001011101111100110011111110010110001011110101111011000010000011001011100111111000011101101000011001101011001110000101111110111110100100100111000110001000000111100001011100010110011010110101011100110100111110001011010100001110110011100110111001101110100100111010101011001000000100101101000001100010000001000010010000110101001111011111101011111110010011001010011000000110110101011011110110111011111111001111001101100101010010011101000010101010011000000011000011000100000101101111100100110011010001111101010001101101010110001010011110101111001100100010101000100111001000011101011111111011100001000110000111010100111101001111000111010010110000111000100111011000100010000010110110111011000111001111000101111011010011100010010111010110100110110110111110110100001110110011001001010010100100011010100111000100111000111100001110000110111010100010010010010101111000110110101111111101011011001110111101111011110011000100011110010010100010001111100110001110000001100100100100101001110001110010000111011110111111111001101010101111000111010011111100100100110100011010011010110101111110011010011110011110000111111001011111000001000010011111100101111010110100000;
    // err_codeword = 1368'b000110110110100000011110100111010110110011001100000010111101100101110100011110111000101110010101111111100001100011000001011100100101110000011101010011110111110010111110110110100101010010011001100001101001010101010110001111001011101111100110011111110010111001011110001011011000010000011001011100111111000011101101000011001101011001110000100111110111110100100100111000110001000000111100001011100010110011010110100001100110100111110001011000100001110010011100110111001101110100100111010101011001000000100101101100001100010010001000010010000100101000111011111111011111110010011001010010000000110110101111011110110111011111111001111001101100101010010011101000010101110011000010011000001010100000101101111100100110011110001111101010001101101010110001010011110101111001100100011101000100111001000011100011111101010100001000110000111110100111101000111000111010110110000111000100111011010100010000010110110111011000111001111000101111011010011100110010101010100100110110110111110110100001111110011001001010010100100011010100111000000111000110100001110000110111010100010010010010101111010110110101110111101011011001110111101111111110000000100011110010010100010001111100110001111000001100100100100101001110001110011000111011110111111111001101010101111000111010011111100100100110100011000011010110101111110011010011110011110000111011001011111000001001010011111100101111010110100000;

    // send_codeword(msg, start_input_enc, data_in_enc);
    // wait (done_enc);
    // receive_codeword(data_out_enc);
    // if (codeword == original) begin
    //   $display("Encoded Successfully");
    // end else begin
    //   $display("Encoder Failure");
    //   $display("%h", codeword);
    //   $display("%h", original);
    // end

    // #20;

    // send_codeword(err_codeword, start_input_dec, data_in_dec);
    // wait (done_dec);
    // receive_codeword(data_out_dec);
    // print_result();
    // #10;

    $display("2: Expected Success");
    // input codeword
    msg = 1368'b001100010111100000101110110011011111100111001010101110001010100011100101000010101110101101110011110101101101011101110010110110011011101110010001100000111010101101000001001101111000000100111100001001100000010011011101101111110110110110000010100100010100100110000110100110010001101001001111001000101001000100000011100101111100011110010010001101010111100011010010010001100010010010000100001100000101101101101110100100010000000111000011010100011010010111101001011010110110001110010001000101011010011001101000110011101000001011010100010100000100111100010001010000000111011010100110101001011101000100011011101000001001110011111010110011000000110001011110100000001000000101101110010001101111100110010010011100110100001100001101000110010111000010000111100110000000111100100001100011001001011001111110100010000001100100011011100101010110001011110100110001100011000011001001000100011010111111011011001111001010100001110010110000000111111101011001110000010001110110100111000110110001011000010001001100111110110010011011001010010010000111;
    original = 1368'b001100010111100000101110110011011111100111001010101110001010100011100101000010101110101101110011110101101101011101110010110110011011101110010001100000111010101101000001001101111000000100111100001001100000010011011101101111110110110110000010100100010100100110000110100110010001101001001111001000101001000100000011100101111100011110010010001101010111100011010010010001100010010010000100001100000101101101101110100100010000000111000011010100011010010111101001011010110110001110010001000101011010011001101000110011101000001011010100010100000100111100010001010000000111011010100110101001011101000100011011101000001001110011111010110011000000110001011110100000001000000101101110010001101111100110010010011100110100001100001101000110010111000010000111100110000000111100100001100011001001011001111110100010000001100100011011100101010110001011110100110001100011000011001001000100011010111111011011001111001010100001110010110000000111111101011001110000010001110110100111000110110001011000010001001100111110110010011011001010010010000111100011011000101000001100011110010001100111011101010010011111000100100110011001010000111010010111110011110101101011000111111011001111001011000110111100111000001110110010101010001101101010010110011100101100111101000101001100101010101100011011110101110100010100000000011000111001111010001101110111011011011100000110010010111110001011100000110000;
    err_codeword = 1368'b001100010111100000101110110011011111100111001010101110001010100011100101000010101010111101110011110101101101011101110010110110011011101110010001100000111010101101000001001101111000000100111101001001100000010011011101101111110110110110001010100100010100100110000110100111010001101001001111001000101001000110000011100101111100011110010010001101010111100011010010010011100010010010000100001100000101101101101110100100010000000111000011010101011010010111101001011010110110001110010010000101011010011001101000110111101000001011010100010101000100111100010001010000010110011010100110101001011101000100011011101000001011110011111010110011000100110011011110100000001000000101101110010011101111100110010010011100110101001100001101000110010111000010000111100110000000111100100011100011001001011001101111100010000001100100011011100001010110001011110100110001100011000011001101000100011010111111011011001111001010100001110010110000000111111101011001110000110001110110100111000111110001011000010001001100111110110010111011001010010010000111100011011000101000001100011110010001100111011101010010011111000100100110010001010000111010010011110011110101101011000111111011001111011111000110111100111000001110110010101010001101101010010110011100101100111101000101001100101010101110011010110101110100010100000000011000111001111010001101110111011011011100000110000010111110001011110000110100;

    send_codeword(msg, start_input_enc, data_in_enc);
    wait (done_enc);
    receive_codeword(data_out_enc);
    if (codeword == original) begin
      $display("Encoded Successfully");
    end else begin
      $display("Encoder Failure");
    end

    #20;

    send_codeword(codeword, start_input_dec, data_in_dec);
    wait (done_dec);
    receive_codeword(data_out_dec);
    print_result();

    #20 $finish;
  end

  task automatic send_codeword;
    input [MAX_CODE_LEN-1:0] codeword;  // Input codeword
    ref start_input;
    ref [MAX_BLOCK_SIZE-1:0] data_in;

    integer i;  // Loop variable
    reg [MAX_BLOCK_SIZE-1:0] temp_num;

    begin
      #10 start_input = 1;
      #10 start_input = 0;
      #10;
      for (i = 0; i < MAX_COLS; i = i + 1) begin
        if (i < cols_in) begin
          temp_num = codeword[MAX_BLOCK_SIZE-1:0];
          temp_num = temp_num << (MAX_BLOCK_SIZE - block_size);
          codeword = codeword >> block_size;
          data_in  = temp_num;
        end else begin
          data_in = 0;
        end
        #10;  // Simulation delay
      end
    end
  endtask

  task automatic receive_codeword;
    ref [MAX_BLOCK_SIZE-1:0] data_out;
    codeword = 0;
    for (i = 0; i < MAX_COLS; i = i + 1) begin
      #10;
      codeword[i*block_size+:MAX_BLOCK_SIZE] = (data_out >> (MAX_BLOCK_SIZE - block_size));
    end
  endtask

  task automatic print_result;
    // Print vectors
    // $display("%h", original);
    // $display("%h", codeword_out);

    if (valid) begin
      $display("\tDecoded output is valid");
      if (codeword == original) begin
        $display("\tCodeword restored");
      end else begin
        $display("\tCodeword not restored");
      end
    end else begin
      $display("\tDecoding failed");
    end
  endtask

endmodule
